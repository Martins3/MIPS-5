
`timescale 1ns / 1ps
module stop_ctrl(
    input clk, 
    input continue,
    input stop
);
endmodule
    