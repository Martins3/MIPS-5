module program_counter(
    input clk, 
    input continue,
    input stop
);
endmodule
    