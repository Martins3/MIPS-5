module stop_ctrl(
    input clk, 
    input continue,
    input stop
);
endmodule
    